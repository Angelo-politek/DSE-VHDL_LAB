LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Es1 IS
PORT ( SW : IN STD_LOGIC_VECTOR(9 DOWNTO 0);
LEDR : OUT STD_LOGIC_VECTOR(9 DOWNTO 0)); 
END Es1;


ARCHITECTURE Behavior OF Es1 IS
BEGIN
LEDR <= SW;
END Behavior;
